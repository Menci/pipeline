`ifndef DECODER_INCLUDED
`define DECODER_INCLUDED

`include "Definitions.sv"
`include "GeneralPurposeRegisters.sv"

`define INST_OP_HIGH        31
`define INST_OP_LOW         26

`define INST_RS_HIGH        25
`define INST_RS_LOW         21
`define INST_RT_HIGH        20
`define INST_RT_LOW         16
`define INST_RD_HIGH        15
`define INST_RD_LOW         11

// R only
`define INST_SH_HIGH      10
`define INST_SH_LOW       6
`define INST_FUNC_HIGH    5
`define INST_FUNC_LOW     0

// I only
`define INST_IMME_HIGH    15
`define INST_IMME_LOW     0

// J only
`define INST_ADDR_HIGH    25
`define INST_ADDR_LOW     0

`define INST_RANGE(inst) `INST_``inst``_HIGH:`INST_``inst``_LOW

typedef enum logic [31:0] {
    ADD     = 32'b000000_????????????????????_100000,
    ADDU    = 32'b000000_????????????????????_100001,
    SUB     = 32'b000000_????????????????????_100010,
    SUBU    = 32'b000000_????????????????????_100011,
    SLL     = 32'b000000_????????????????????_000000,
    SRL     = 32'b000000_????????????????????_000010,
    SRA     = 32'b000000_????????????????????_000011,
    SLLV    = 32'b000000_????????????????????_000100,
    SRLV    = 32'b000000_????????????????????_000110,
    SRAV    = 32'b000000_????????????????????_000111,
    AND     = 32'b000000_????????????????????_100100,
    OR      = 32'b000000_????????????????????_100101,
    XOR     = 32'b000000_????????????????????_100110,
    NOR     = 32'b000000_????????????????????_100111,
    SLT     = 32'b000000_????????????????????_101010,
    SLTU    = 32'b000000_????????????????????_101011,

    ADDI    = 32'b001000_????????????????????_??????,
    ADDIU   = 32'b001001_????????????????????_??????,
    ANDI    = 32'b001100_????????????????????_??????,
    ORI     = 32'b001101_????????????????????_??????,
    XORI    = 32'b001110_????????????????????_??????,
    SLTI    = 32'b001010_????????????????????_??????,
    SLTIU   = 32'b001011_????????????????????_??????,

    LUI     = 32'b001111_????????????????????_??????,

    MULT    = 32'b000000_????????????????????_011000,
    MULTU   = 32'b000000_????????????????????_011001,
    DIV     = 32'b000000_????????????????????_011010,
    DIVU    = 32'b000000_????????????????????_011011,
    MFHI    = 32'b000000_????????????????????_010000,
    MTHI    = 32'b000000_????????????????????_010001,
    MFLO    = 32'b000000_????????????????????_010010,
    MTLO    = 32'b000000_????????????????????_010011,

    BEQ     = 32'b000100_????????????????????_??????,
    BNE     = 32'b000101_????????????????????_??????,
    BLEZ    = 32'b000110_????????????????????_??????,
    BGTZ    = 32'b000111_????????????????????_??????,
    BGEZ    = 32'b000001_?????00001??????????_??????,
    BLTZ    = 32'b000001_?????00000??????????_??????,

    JR      = 32'b000000_????????????????????_001000,
    JALR    = 32'b000000_????????????????????_001001,
    J       = 32'b000010_????????????????????_??????,
    JAL     = 32'b000011_????????????????????_??????,

    LB      = 32'b100000_????????????????????_??????,
    LBU     = 32'b100100_????????????????????_??????,
    LH      = 32'b100001_????????????????????_??????,
    LHU     = 32'b100101_????????????????????_??????,
    LW      = 32'b100011_????????????????????_??????,
    SB      = 32'b101000_????????????????????_??????,
    SH      = 32'b101001_????????????????????_??????,
    SW      = 32'b101011_????????????????????_??????,

    SYSCALL = 32'b000000_????????????????????_001100
} instruction_code_t;

typedef logic [`INST_SH_HIGH - `INST_SH_LOW:0] shift_amount_t;
typedef logic [`INST_IMME_HIGH - `INST_IMME_LOW:0] immediate_t;
typedef logic [`INST_ADDR_HIGH - `INST_ADDR_LOW:0] absolute_jump_input_t;

typedef struct packed {
    instruction_code_t instructionCode;
    register_id_t registerS;
    register_id_t registerT;
    register_id_t registerD;
    shift_amount_t shiftAmount;
    immediate_t immediate;
    absolute_jump_input_t absoluteJumpInput;
} instruction_t;

// Include the file after enum
`include "Debug.sv"

function instruction_t parseInstruction(int_t instructionData);
    instruction_t instruction;

`ifndef DEBUG_INSTRUCTION_CODE_ENUM
    instruction.instructionCode = instruction_code_t'(instructionData);
`else
    instruction.instructionCode = getInstructionCode(instructionData);
`endif
    instruction.registerS = register_id_t'(instructionData[`INST_RANGE(RS)]);
    instruction.registerT = register_id_t'(instructionData[`INST_RANGE(RT)]);
    instruction.registerD = register_id_t'(instructionData[`INST_RANGE(RD)]);
    instruction.shiftAmount = instructionData[`INST_RANGE(SH)];
    instruction.immediate = instructionData[`INST_RANGE(IMME)];
    instruction.absoluteJumpInput = instructionData[`INST_RANGE(ADDR)];

    return instruction;
endfunction

`endif // DECODER_INCLUDED
